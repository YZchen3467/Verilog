/*Getting Started*/
module top_module( output one );

// Insert your code here
    assign one = 1;

endmodule

///////////////////////////////////

/*Output Zero*/
module top_module(output zero)

	assign zero = 0;

endmodule